`timescale 1ps/1ps

module InstructionMemory(
    input PCF,
    output logic InstrF
);
endmodule