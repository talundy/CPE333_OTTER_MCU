`timescale 1ps/1ps

module PC(
    input CLK,
    input PCFPrime,
    output logic PCF
);
endmodule