`timescale 1ps/1ps

module AddFour(
    input PCF,
    output logic PCPlusFour
); 
endmodule