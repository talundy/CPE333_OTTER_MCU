`timescale 1ps/1ps

module PCMux (
    input PCSourceE,        // enable signal from E stage 
    input PCPlus4F,         
    input PCTargetE,        
    output logic PCFPrime
);
endmodule